/* A simple AND gate File: and2.v */
module andgate(y,a,b,);
input a,b;
output y;
assign y=a&b;
endmodule
