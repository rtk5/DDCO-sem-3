module andgate (y,a, );  
input a;
output y;
assign y = !a;
endmodule
